`timescale 1ns/1ns
//`include "fsm.v"
module stimulus_2;
reg clk;
//reg rst1;
reg rst;
reg [15:0] x;
wire z;

wire try;

wire reset_try;
fsm UUT(clk,rst,x,z,try,reset_try);

initial
  begin
    $dumpfile("stimulus_tb3.vcd");
    $dumpvars;
  end


initial
    clk=1'b0;
always
    #5 clk =~clk;
initial
begin
    rst=1'b1;
    x=16'b1111111111111111;
    #10 rst=1'b0;
    #10 x=16'b1101111101101111;
    #10 x=16'b1101111101101111;
    #10 x=16'b1101111101101111;
    #10 x=16'b1101111101101111;
    #10 rst=1'b0;	
    #10 x=16'b1101111101101111;
    #10 x=16'b1111110110101111;
    #10 x=16'b1101011011111111;
    #10 x=16'b0000000000000000;
    #10 x=16'b1111011011011011;
    #10 x=16'b1111110110101111;
    #10 x=16'b1101011011111111;
    #10 x=16'b1111011011011011;
    #10 x=16'b1010101010101010;
    #10 x=16'b0101010101010101;
    #10 x=16'b1100110011001100;
    #10 x=16'b0011001100110011;	
    #10 x=16'b0000000000000000;
    #10 x=16'b1000000000000000;
    rst=1'b1;
    x=16'b1111111111111111;
    #10 rst=1'b0;
    #10 x=16'b0000000000000000;
    #10 x=16'b0000000000000000;
    #10 x=16'b0000000000000000;
    #10 x=16'b0000000000000000;
    #10 x=16'b0000000000000000;
    #10 x=16'b0000000000000000;
    #10 x=16'b1111111111111110;
    #10 x=16'b1111011111111111;
    rst=1'b1;
    #10 x=16'b1101101111111111;
    #10 x=16'b1101111101101111;
    rst=1'b0;
    #10 x=16'b0000000000000000;
    #10 x=16'b0000000000000000;
    #10 x=16'b0000000000000000;
    #10 x=16'b0000000000000000;
    #10 x=16'b0000000000000000;
    #10 x=16'b0000000000000000;
    #10 x=16'b1101111101101111;
    #10 x=16'b1101111101101111;
    #10 x=16'b1101111101101111;
    #10 x=16'b1101111101101111;
    #10 x=16'b1111110110101111;
    #10 x=16'b1101011011111111;
    #10 x=16'b1111011011011011;
    #10 x=16'b1111110110101111;
    #10 x=16'b1101011011111111;
    #10 x=16'b1111011011011011;
    #10 x=16'b0000000000000000;
    #20 $finish;
end
initial
    $monitor($time," Output z= %d and input x=%d and try=%d and reset_try=%d",z,x,try,reset_try);
endmodule
